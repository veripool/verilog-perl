// DESCRIPTION: Verilog-Perl: Example Verilog for testing package
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2000-2012 by Wilson Snyder.

`ifndef V_HIER_INC_VH
`define V_HIER_INC_VH  // Guard

`define hsub v_hier_sub

`endif  // Guard
