// DESCRIPTION: Verilog::Preproc: Example source code
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2012-2012 by Wilson Snyder.
//
// Test -F option in vppreproc.

module bar(output wire y, input wire x);
   assign y = x;
endmodule // bar
