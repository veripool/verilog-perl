// DESCRIPTION: Verilog::Preproc: Example source code
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2000-2010 by Wilson Snyder.

module t_86_vhier_tick;

   `define t_86_vhier_tick_sub FOOBAR_NOT_FOUND
   t_86_vhier_tick_sub sub ();

endmodule
